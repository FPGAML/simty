library ieee;
use ieee.std_logic_1164.all;

entity Instruction_ROM is
	port (
		clock : in std_logic;
		addr : in std_logic_vector(7 downto 0);
		data : out std_logic_vector(31 downto 0)
	);
end entity;

architecture structural of Instruction_ROM is
	signal addr_1 : std_logic_vector(7 downto 0);
begin
	process(clock)
	begin
		if rising_edge(clock) then
			case addr is
				when X"00" => data <= X"464c457f";
				when X"01" => data <= X"00010101";
				when X"02" => data <= X"00000000";
				when X"03" => data <= X"00000000";
				when X"04" => data <= X"00f30002";
				when X"05" => data <= X"00000001";
				when X"06" => data <= X"00000200";
				when X"07" => data <= X"00000034";
				when X"08" => data <= X"0000033c";
				when X"09" => data <= X"00000000";
				when X"0a" => data <= X"00200034";
				when X"0b" => data <= X"00280001";
				when X"0c" => data <= X"00020005";
				when X"0d" => data <= X"00000001";
				when X"0e" => data <= X"00000000";
				when X"0f" => data <= X"00000000";
				when X"10" => data <= X"00000000";
				when X"11" => data <= X"00000234";
				when X"12" => data <= X"00000234";
				when X"13" => data <= X"00000005";
				when X"14" => data <= X"00001000";
				when X"15" => data <= X"00000000";
				when X"16" => data <= X"00000000";
				when X"17" => data <= X"00000000";
				when X"18" => data <= X"00000000";
				when X"19" => data <= X"00000000";
				when X"1a" => data <= X"00000000";
				when X"1b" => data <= X"00000000";
				when X"1c" => data <= X"00000000";
				when X"1d" => data <= X"00000000";
				when X"1e" => data <= X"00000000";
				when X"1f" => data <= X"00000000";
				when X"20" => data <= X"00000000";
				when X"21" => data <= X"00000000";
				when X"22" => data <= X"00000000";
				when X"23" => data <= X"00000000";
				when X"24" => data <= X"00000000";
				when X"25" => data <= X"00000000";
				when X"26" => data <= X"00000000";
				when X"27" => data <= X"00000000";
				when X"28" => data <= X"00000000";
				when X"29" => data <= X"00000000";
				when X"2a" => data <= X"00000000";
				when X"2b" => data <= X"00000000";
				when X"2c" => data <= X"00000000";
				when X"2d" => data <= X"00000000";
				when X"2e" => data <= X"00000000";
				when X"2f" => data <= X"00000000";
				when X"30" => data <= X"00000000";
				when X"31" => data <= X"00000000";
				when X"32" => data <= X"00000000";
				when X"33" => data <= X"00000000";
				when X"34" => data <= X"00000000";
				when X"35" => data <= X"00000000";
				when X"36" => data <= X"00000000";
				when X"37" => data <= X"00000000";
				when X"38" => data <= X"00000000";
				when X"39" => data <= X"00000000";
				when X"3a" => data <= X"00000000";
				when X"3b" => data <= X"00000000";
				when X"3c" => data <= X"00000000";
				when X"3d" => data <= X"00000000";
				when X"3e" => data <= X"00000000";
				when X"3f" => data <= X"00000000";
				when X"40" => data <= X"00000000";
				when X"41" => data <= X"00000000";
				when X"42" => data <= X"00000000";
				when X"43" => data <= X"00000000";
				when X"44" => data <= X"00000000";
				when X"45" => data <= X"00000000";
				when X"46" => data <= X"00000000";
				when X"47" => data <= X"00000000";
				when X"48" => data <= X"00000000";
				when X"49" => data <= X"00000000";
				when X"4a" => data <= X"00000000";
				when X"4b" => data <= X"00000000";
				when X"4c" => data <= X"00000000";
				when X"4d" => data <= X"00000000";
				when X"4e" => data <= X"00000000";
				when X"4f" => data <= X"00000000";
				when X"50" => data <= X"00000000";
				when X"51" => data <= X"00000000";
				when X"52" => data <= X"00000000";
				when X"53" => data <= X"00000000";
				when X"54" => data <= X"00000000";
				when X"55" => data <= X"00000000";
				when X"56" => data <= X"00000000";
				when X"57" => data <= X"00000000";
				when X"58" => data <= X"00000000";
				when X"59" => data <= X"00000000";
				when X"5a" => data <= X"00000000";
				when X"5b" => data <= X"00000000";
				when X"5c" => data <= X"00000000";
				when X"5d" => data <= X"00000000";
				when X"5e" => data <= X"00000000";
				when X"5f" => data <= X"00000000";
				when X"60" => data <= X"00000000";
				when X"61" => data <= X"00000000";
				when X"62" => data <= X"00000000";
				when X"63" => data <= X"00000000";
				when X"64" => data <= X"00000000";
				when X"65" => data <= X"00000000";
				when X"66" => data <= X"00000000";
				when X"67" => data <= X"00000000";
				when X"68" => data <= X"00000000";
				when X"69" => data <= X"00000000";
				when X"6a" => data <= X"00000000";
				when X"6b" => data <= X"00000000";
				when X"6c" => data <= X"00000000";
				when X"6d" => data <= X"00000000";
				when X"6e" => data <= X"00000000";
				when X"6f" => data <= X"00000000";
				when X"70" => data <= X"00000000";
				when X"71" => data <= X"00000000";
				when X"72" => data <= X"00000000";
				when X"73" => data <= X"00000000";
				when X"74" => data <= X"00000000";
				when X"75" => data <= X"00000000";
				when X"76" => data <= X"00000000";
				when X"77" => data <= X"00000000";
				when X"78" => data <= X"00000000";
				when X"79" => data <= X"00000000";
				when X"7a" => data <= X"00000000";
				when X"7b" => data <= X"00000000";
				when X"7c" => data <= X"00000000";
				when X"7d" => data <= X"00000000";
				when X"7e" => data <= X"00000000";
				when X"7f" => data <= X"00000000";
				when X"80" => data <= X"02a00613";
				when X"81" => data <= X"01010437";
				when X"82" => data <= X"10140413";
				when X"83" => data <= X"000014b7";
				when X"84" => data <= X"00000537";
				when X"85" => data <= X"f10025f3";
				when X"86" => data <= X"00259593";
				when X"87" => data <= X"00b502b3";
				when X"88" => data <= X"00c2a023";
				when X"89" => data <= X"02058593";
				when X"8a" => data <= X"fe95cae3";
				when X"8b" => data <= X"00860633";
				when X"8c" => data <= X"fe5ff06f";
				when X"8d" => data <= X"00000000";
				when X"8e" => data <= X"00000000";
				when X"8f" => data <= X"00000000";
				when X"90" => data <= X"00000000";
				when X"91" => data <= X"00000000";
				when X"92" => data <= X"00000000";
				when X"93" => data <= X"00000000";
				when X"94" => data <= X"00000000";
				when X"95" => data <= X"00000000";
				when X"96" => data <= X"00000000";
				when X"97" => data <= X"00000000";
				when X"98" => data <= X"00000000";
				when X"99" => data <= X"00000000";
				when X"9a" => data <= X"00000000";
				when X"9b" => data <= X"00000000";
				when X"9c" => data <= X"00000000";
				when X"9d" => data <= X"00000000";
				when X"9e" => data <= X"00000000";
				when X"9f" => data <= X"00000000";
				when X"a0" => data <= X"00000000";
				when X"a1" => data <= X"00000000";
				when X"a2" => data <= X"00000000";
				when X"a3" => data <= X"00000000";
				when X"a4" => data <= X"00000000";
				when X"a5" => data <= X"00000000";
				when X"a6" => data <= X"00000000";
				when X"a7" => data <= X"00000000";
				when X"a8" => data <= X"00000000";
				when X"a9" => data <= X"00000000";
				when X"aa" => data <= X"00000000";
				when X"ab" => data <= X"00000000";
				when X"ac" => data <= X"00000000";
				when X"ad" => data <= X"00000000";
				when X"ae" => data <= X"00000000";
				when X"af" => data <= X"00000000";
				when X"b0" => data <= X"00000000";
				when X"b1" => data <= X"00000000";
				when X"b2" => data <= X"00000000";
				when X"b3" => data <= X"00000000";
				when X"b4" => data <= X"00000000";
				when X"b5" => data <= X"00000000";
				when X"b6" => data <= X"00000000";
				when X"b7" => data <= X"00000000";
				when X"b8" => data <= X"00000000";
				when X"b9" => data <= X"00000000";
				when X"ba" => data <= X"00000000";
				when X"bb" => data <= X"00000000";
				when X"bc" => data <= X"00000000";
				when X"bd" => data <= X"00000000";
				when X"be" => data <= X"00000000";
				when X"bf" => data <= X"00000000";
				when X"c0" => data <= X"00000000";
				when X"c1" => data <= X"00000000";
				when X"c2" => data <= X"00000000";
				when X"c3" => data <= X"00000000";
				when X"c4" => data <= X"00000000";
				when X"c5" => data <= X"00000000";
				when X"c6" => data <= X"00000000";
				when X"c7" => data <= X"00000000";
				when X"c8" => data <= X"00000000";
				when X"c9" => data <= X"00000000";
				when X"ca" => data <= X"00000000";
				when X"cb" => data <= X"00000000";
				when X"cc" => data <= X"00000000";
				when X"cd" => data <= X"00000000";
				when X"ce" => data <= X"00000000";
				when X"cf" => data <= X"00000000";
				when X"d0" => data <= X"00000000";
				when X"d1" => data <= X"00000000";
				when X"d2" => data <= X"00000000";
				when X"d3" => data <= X"00000000";
				when X"d4" => data <= X"00000000";
				when X"d5" => data <= X"00000000";
				when X"d6" => data <= X"00000000";
				when X"d7" => data <= X"00000000";
				when X"d8" => data <= X"00000000";
				when X"d9" => data <= X"00000000";
				when X"da" => data <= X"00000000";
				when X"db" => data <= X"00000000";
				when X"dc" => data <= X"00000000";
				when X"dd" => data <= X"00000000";
				when X"de" => data <= X"00000000";
				when X"df" => data <= X"00000000";
				when X"e0" => data <= X"00000000";
				when X"e1" => data <= X"00000000";
				when X"e2" => data <= X"00000000";
				when X"e3" => data <= X"00000000";
				when X"e4" => data <= X"00000000";
				when X"e5" => data <= X"00000000";
				when X"e6" => data <= X"00000000";
				when X"e7" => data <= X"00000000";
				when X"e8" => data <= X"00000000";
				when X"e9" => data <= X"00000000";
				when X"ea" => data <= X"00000000";
				when X"eb" => data <= X"00000000";
				when X"ec" => data <= X"00000000";
				when X"ed" => data <= X"00000000";
				when X"ee" => data <= X"00000000";
				when X"ef" => data <= X"00000000";
				when X"f0" => data <= X"00000000";
				when X"f1" => data <= X"00000000";
				when X"f2" => data <= X"00000000";
				when X"f3" => data <= X"00000000";
				when X"f4" => data <= X"00000000";
				when X"f5" => data <= X"00000000";
				when X"f6" => data <= X"00000000";
				when X"f7" => data <= X"00000000";
				when X"f8" => data <= X"00000000";
				when X"f9" => data <= X"00000000";
				when X"fa" => data <= X"00000000";
				when X"fb" => data <= X"00000000";
				when X"fc" => data <= X"00000000";
				when X"fd" => data <= X"00000000";
				when X"fe" => data <= X"00000000";
				when X"ff" => data <= X"00000000";
				when others => data <= (others => '-');
			end case;
		end if;
	end process;
end architecture;
